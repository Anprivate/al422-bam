library verilog;
use verilog.vl_types.all;
entity al422_bam_vlg_tst is
end al422_bam_vlg_tst;
